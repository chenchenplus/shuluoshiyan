module ALUController(input [5:0]OpCode,
           input [5:0] Funct,
           output reg [4:0] ALUCtrl,
           output reg Sign
);
always @(*) begin
    case(OpCode)
    6'h00:begin
         case(Funct)
         //add
         6'h20:begin
               ALUCtrl=5'b00000;
               Sign=1'b1;
               end
         //addu
         6'h21:begin
               ALUCtrl=5'b00000;
               Sign=1'b0;
               end
         //sub
         6'h22:begin
               ALUCtrl=5'b00001;
               Sign=1'b1;
               end
         //subu
         6'h23:begin
               ALUCtrl=5'b00001;
               Sign=1'b0;
               end
         //and
         6'h24:begin
               ALUCtrl=5'b00010;
               Sign=1'b1;
               end
         //or
         6'h25:begin
               ALUCtrl=5'b00011;
               Sign=1'b1;
               end
         //xor
         6'h26:begin
               ALUCtrl=5'b00100;
               Sign=1'b1;
               end
         //nor
         6'h27:begin
               ALUCtrl=5'b00101;
               Sign=1'b1;
               end
         //sll
         6'h00:begin
               ALUCtrl=5'b00110;
               Sign=1'b0;
               end
         //srl
         6'h02:begin
               ALUCtrl=5'b00111;
               Sign=1'b0;
               end
         //sra
         6'h03:begin
               ALUCtrl=5'b01000;
               Sign=1'b1;
               end
         //slt
         6'h2a:begin
               ALUCtrl=5'b01001;
               Sign=1'b1;
               end
         //sltu
         6'h2b:begin
               ALUCtrl=5'b01001;
               Sign=1'b0;
               end
         endcase
         end
    //lw
    6'h23:begin
          ALUCtrl=5'b00000;
          Sign=1'b1;
          end
    //sw
    6'h2b:begin
          ALUCtrl=5'b00000;
          Sign=1'b1;
          end
    //addi
    6'h08:begin
          ALUCtrl=5'b00000;
          Sign=1'b1;
          end
    //addiu
    6'h09:begin
          ALUCtrl=5'b00000;
          Sign=1'b0;
          end
    //andi
    6'h0c:begin
          ALUCtrl=5'b00010;
          Sign=1'b0;
          end
    //slti
    6'h0a:begin
          ALUCtrl=5'b01001;
          Sign=1'b1;
          end
    //sltiu
    6'h0b:begin
          ALUCtrl=5'b01001;
          Sign=1'b0;
          end
    //beq
    6'h04:begin
          ALUCtrl=5'b00001;
          Sign=1'b1;
          end
    endcase
end
endmodule